module example_block
#(
    parameter PARAM    = 1,
              FOO            = 2,
              BARFLUG                = 4,
              G                      = 5
)
    (// I/O
     input     reset_n,
     input     clk,
     input     a, b,
     output reg c
    );
endmodule

